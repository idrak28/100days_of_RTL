library verilog;
use verilog.vl_types.all;
entity seq_TB is
end seq_TB;
