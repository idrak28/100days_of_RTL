library verilog;
use verilog.vl_types.all;
entity lab2tb is
end lab2tb;
