library verilog;
use verilog.vl_types.all;
entity lab2 is
    port(
        i               : in     vl_logic;
        clk             : in     vl_logic;
        \out\           : out    vl_logic
    );
end lab2;
